module megavliw #(
    parameter VLIW_WIDTH = 128,
) (
    input wire clk,
    input wire rst
);
endmodule